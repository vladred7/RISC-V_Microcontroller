module cpu_top #(
    parameter ADDR_WIDTH = 5,
    parameter DATA_WIDTH = 32
)(
	input clk,    // Clock
	
);

   import pkg_cpu_typedefs::*;

endmodule : cpu_top