module cpu_fsm_decoder (
	input clk,    // Clock
	input clk_en, // Clock Enable
	input rst_n,  // Asynchronous reset active low
	
);
   
   import pkg_cpu_typedefs::*;

endmodule : cpu_fsm_decoder