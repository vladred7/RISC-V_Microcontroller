module sfr_map #(
   parameter SFR_WIDTH              = 32
)(
   //    Input ports definition
   input                   sys_clk,
   input                   sys_clk_en,
   input                   sys_rst_n
   //input                   sfr_wen,
   //input  [SFR_WIDTH-1:0]  sfr_din,
   //    Output ports definition
   //output [SFR_WIDTH-1:0]  sfr_dout,
   //output [SFR_WIDTH-1:0]  sfr_rdonly_dout
);

endmodule : sfr_map